module num_switch (
    input [3:0] digit,
    input [4:0]y,
    input [4:0]x,
    output reg has_color
);
reg [19:0] num_line;
always @(*) begin
        case (digit)
            4'b0000:
            begin
                case (y)
                     0: num_line=20'b00000000000000000000;
                     1: num_line=20'b00000000000000000000;
                     2: num_line=20'b00000000000000000000;
                     3: num_line=20'b00000000000000000000;
                     4: num_line=20'b00000000000000000000;
                     5: num_line=20'b00000000000000000000;
                     6: num_line=20'b00000000000000000000;
                     7: num_line=20'b00000000000000000000;
                     8: num_line=20'b00000000000000000000;
                     9: num_line=20'b00001100000000000000;
                    10: num_line=20'b00011100000000000000;
                    11: num_line=20'b00111111000000000000;
                    12: num_line=20'b01111111000000000000;
                    13: num_line=20'b01111111000000000000;
                    14: num_line=20'b01110111100000000000;
                    15: num_line=20'b11100011100000000000;
                    16: num_line=20'b11100011100000000000;
                    17: num_line=20'b11100011100000000000;
                    18: num_line=20'b11100011100000000000;
                    19: num_line=20'b11100001100000000000;
                    20: num_line=20'b11100001100000000000;
                    21: num_line=20'b11100001100000000000;
                    22: num_line=20'b11100001100000000000;
                    23: num_line=20'b11100001100000000000;
                    24: num_line=20'b11100011100000000000;
                    25: num_line=20'b11100011100000000000;
                    26: num_line=20'b11100011100000000000;
                    27: num_line=20'b11110011100000000000;
                    28: num_line=20'b01110111100000000000;
                    29: num_line=20'b01110111100000000000;
                    30: num_line=20'b01111111000000000000;
                    31: num_line=20'b00111110000000000000;
                    default: num_line=20'b00000000000000000000;
                endcase
            end
            4'b0001: //1
            begin
                case (y)
                     0: num_line=20'b00000000000000000000;
                     1: num_line=20'b00000000000000000000;
                     2: num_line=20'b00000000000000000000;
                     3: num_line=20'b00000000000000000000;
                     4: num_line=20'b00000000000000000000;
                     5: num_line=20'b00000000000000000000;
                     6: num_line=20'b00000000000000000000;
                     7: num_line=20'b00000000000000000000;
                     8: num_line=20'b00000000000000000000;
                     9: num_line=20'b00001100000000000000;
                    10: num_line=20'b00001100000000000000;
                    11: num_line=20'b00011100000000000000;
                    12: num_line=20'b00111100000000000000;
                    13: num_line=20'b00111100000000000000;
                    14: num_line=20'b01111100000000000000;
                    15: num_line=20'b01111100000000000000;
                    16: num_line=20'b01111100000000000000;
                    17: num_line=20'b01111100000000000000;
                    18: num_line=20'b00011100000000000000;
                    19: num_line=20'b00011100000000000000;
                    20: num_line=20'b00011100000000000000;
                    21: num_line=20'b00011100000000000000;
                    22: num_line=20'b00011100000000000000;
                    23: num_line=20'b00011100000000000000;
                    24: num_line=20'b00011100000000000000;
                    25: num_line=20'b00011100000000000000;
                    26: num_line=20'b00011100000000000000;
                    27: num_line=20'b00011100000000000000;
                    28: num_line=20'b00011110000000000000;
                    29: num_line=20'b00011110000000000000;
                    30: num_line=20'b00111111000000000000;
                    31: num_line=20'b00111111000000000000;
                    default: num_line=20'b00000000000000000000;
                endcase
            end
            4'b0010: begin //2
                case (y)
                     0: num_line=20'b00000000000000000000;
                     1: num_line=20'b00000000000000000000;
                     2: num_line=20'b00000000000000000000;
                     3: num_line=20'b00000000000000000000;
                     4: num_line=20'b00000000000000000000;
                     5: num_line=20'b00000000000000000000;
                     6: num_line=20'b00000000000000000000;
                     7: num_line=20'b00000000000000000000;
                     8: num_line=20'b00000000000000000000;
                     9: num_line=20'b00011100000000000000;
                    10: num_line=20'b00011110000000000000;
                    11: num_line=20'b00111111000000000000;
                    12: num_line=20'b01111111100000000000;
                    13: num_line=20'b01111111100000000000;
                    14: num_line=20'b01111111100000000000;
                    15: num_line=20'b11100011100000000000;
                    16: num_line=20'b11100011100000000000;
                    17: num_line=20'b11100011100000000000;
                    18: num_line=20'b00000011100000000000;
                    19: num_line=20'b00000111100000000000;
                    20: num_line=20'b00001111100000000000;
                    21: num_line=20'b00001111000000000000;
                    22: num_line=20'b00001111000000000000;
                    23: num_line=20'b00011110000000000000;
                    24: num_line=20'b00011110000000000000;
                    25: num_line=20'b00111100100000000000;
                    26: num_line=20'b00111000100000000000;
                    27: num_line=20'b01111001100000000000;
                    28: num_line=20'b11111111100000000000;
                    29: num_line=20'b11111111100000000000;
                    30: num_line=20'b11111111100000000000;
                    31: num_line=20'b11111111100000000000;
                    default: num_line=20'b00000000000000000000;
                endcase
            end
            4'b0011:begin
                case (y)
                     0: num_line=20'b00000000000000000000;
                     1: num_line=20'b00000000000000000000;
                     2: num_line=20'b00000000000000000000;
                     3: num_line=20'b00000000000000000000;
                     4: num_line=20'b00000000000000000000;
                     5: num_line=20'b00000000000000000000;
                     6: num_line=20'b00000000000000000000;
                     7: num_line=20'b00000000000000000000;
                     8: num_line=20'b00000000000000000000;
                     9: num_line=20'b00001110000000000000;
                    10: num_line=20'b00001110000000000000;
                    11: num_line=20'b00111111000000000000;
                    12: num_line=20'b01111111000000000000;
                    13: num_line=20'b01111111000000000000;
                    14: num_line=20'b01111111000000000000;
                    15: num_line=20'b01100111000000000000;
                    16: num_line=20'b01100111000000000000;
                    17: num_line=20'b01001111000000000000;
                    18: num_line=20'b00001110000000000000;
                    19: num_line=20'b00011111100000000000;
                    20: num_line=20'b00011111100000000000;
                    21: num_line=20'b00011111100000000000;
                    22: num_line=20'b00011111100000000000;
                    23: num_line=20'b00000011100000000000;
                    24: num_line=20'b00000011100000000000;
                    25: num_line=20'b00000011100000000000;
                    26: num_line=20'b00000011100000000000;
                    27: num_line=20'b00000011100000000000;
                    28: num_line=20'b11110111100000000000;
                    29: num_line=20'b11110111100000000000;
                    30: num_line=20'b11111111000000000000;
                    31: num_line=20'b11111110000000000000;
                    default: num_line=20'b00000000000000000000;
                endcase
            end 
            4'b0100: begin
                case (y)
                     0: num_line=20'b00000000000000000000;
                     1: num_line=20'b00000000000000000000;
                     2: num_line=20'b00000000000000000000;
                     3: num_line=20'b00000000000000000000;
                     4: num_line=20'b00000000000000000000;
                     5: num_line=20'b00000000000000000000;
                     6: num_line=20'b00000000000000000000;
                     7: num_line=20'b00000000000000000000;
                     8: num_line=20'b00000000000000000000;
                     9: num_line=20'b00000011000000000000;
                    10: num_line=20'b00000011000000000000;
                    11: num_line=20'b00000111000000000000;
                    12: num_line=20'b00001111000000000000;
                    13: num_line=20'b00001111000000000000;
                    14: num_line=20'b00001111000000000000;
                    15: num_line=20'b00011111000000000000;
                    16: num_line=20'b00011111000000000000;
                    17: num_line=20'b00111111000000000000;
                    18: num_line=20'b00111111000000000000;
                    19: num_line=20'b00111111000000000000;
                    20: num_line=20'b01110111000000000000;
                    21: num_line=20'b01110111000000000000;
                    22: num_line=20'b11110111000000000000;
                    23: num_line=20'b11111111110000000000;
                    24: num_line=20'b11111111110000000000;
                    25: num_line=20'b11111111110000000000;
                    26: num_line=20'b11111111110000000000;
                    27: num_line=20'b11111111110000000000;
                    28: num_line=20'b00000111000000000000;
                    29: num_line=20'b00000111000000000000;
                    30: num_line=20'b00000111000000000000;
                    31: num_line=20'b00000111000000000000;
                    default: num_line=20'b00000000000000000000;
                endcase
            end
            4'b0101: begin
                case (y)
                     0: num_line=20'b00000000000000000000;
                     1: num_line=20'b00000000000000000000;
                     2: num_line=20'b00000000000000000000;
                     3: num_line=20'b00000000000000000000;
                     4: num_line=20'b00000000000000000000;
                     5: num_line=20'b00000000000000000000;
                     6: num_line=20'b00000000000000000000;
                     7: num_line=20'b00000000000000000000;
                     8: num_line=20'b00000000000000000000;
                     9: num_line=20'b00111111000000000000;
                    10: num_line=20'b00111111000000000000;
                    11: num_line=20'b00111111000000000000;
                    12: num_line=20'b00111111000000000000;
                    13: num_line=20'b00111111000000000000;
                    14: num_line=20'b00111111000000000000;
                    15: num_line=20'b00110000000000000000;
                    16: num_line=20'b00110000000000000000;
                    17: num_line=20'b00111110000000000000;
                    18: num_line=20'b00111110000000000000;
                    19: num_line=20'b00111111000000000000;
                    20: num_line=20'b00111111100000000000;
                    21: num_line=20'b00111111100000000000;
                    22: num_line=20'b00111111100000000000;
                    23: num_line=20'b00000011100000000000;
                    24: num_line=20'b00000011100000000000;
                    25: num_line=20'b00000011100000000000;
                    26: num_line=20'b00000011100000000000;
                    27: num_line=20'b00000011100000000000;
                    28: num_line=20'b01110111100000000000;
                    29: num_line=20'b01110111100000000000;
                    30: num_line=20'b01111111000000000000;
                    31: num_line=20'b01111111000000000000;
                    default: num_line=20'b00000000000000000000;
                endcase
            end
            4'b0110:begin
                case (y)
                     0: num_line=20'b00000000000000000000;
                     1: num_line=20'b00000000000000000000;
                     2: num_line=20'b00000000000000000000;
                     3: num_line=20'b00000000000000000000;
                     4: num_line=20'b00000000000000000000;
                     5: num_line=20'b00000000000000000000;
                     6: num_line=20'b00000000000000000000;
                     7: num_line=20'b00000000000000000000;
                     8: num_line=20'b00000000000000000000;
                     9: num_line=20'b00000001000000000000;
                    10: num_line=20'b00000011000000000000;
                    11: num_line=20'b00001111000000000000;
                    12: num_line=20'b00011111000000000000;
                    13: num_line=20'b00011111000000000000;
                    14: num_line=20'b00111110000000000000;
                    15: num_line=20'b00111100000000000000;
                    16: num_line=20'b01111100000000000000;
                    17: num_line=20'b01111000000000000000;
                    18: num_line=20'b01110000000000000000;
                    19: num_line=20'b01111111000000000000;
                    20: num_line=20'b11111111100000000000;
                    21: num_line=20'b11111111100000000000;
                    22: num_line=20'b11101111100000000000;
                    23: num_line=20'b11100011100000000000;
                    24: num_line=20'b11100011100000000000;
                    25: num_line=20'b11100011100000000000;
                    26: num_line=20'b11100011100000000000;
                    27: num_line=20'b11110011100000000000;
                    28: num_line=20'b01110111100000000000;
                    29: num_line=20'b01110111100000000000;
                    30: num_line=20'b01111111100000000000;
                    31: num_line=20'b00111111000000000000;
                    default: num_line=20'b00000000000000000000;
                endcase
            end 
            4'b0111: begin
                case (y)
                     0: num_line=20'b00000000000000000000;
                     1: num_line=20'b00000000000000000000;
                     2: num_line=20'b00000000000000000000;
                     3: num_line=20'b00000000000000000000;
                     4: num_line=20'b00000000000000000000;
                     5: num_line=20'b00000000000000000000;
                     6: num_line=20'b00000000000000000000;
                     7: num_line=20'b00000000000000000000;
                     8: num_line=20'b00000000000000000000;
                     9: num_line=20'b01111111100000000000;
                    10: num_line=20'b11111111100000000000;
                    11: num_line=20'b11111111100000000000;
                    12: num_line=20'b11111111100000000000;
                    13: num_line=20'b11111111100000000000;
                    14: num_line=20'b11111111100000000000;
                    15: num_line=20'b11000011100000000000;
                    16: num_line=20'b11000011100000000000;
                    17: num_line=20'b00000111000000000000;
                    18: num_line=20'b00000111000000000000;
                    19: num_line=20'b00000111000000000000;
                    20: num_line=20'b00000110000000000000;
                    21: num_line=20'b00000110000000000000;
                    22: num_line=20'b00001110000000000000;
                    23: num_line=20'b00001110000000000000;
                    24: num_line=20'b00001110000000000000;
                    25: num_line=20'b00001100000000000000;
                    26: num_line=20'b00001100000000000000;
                    27: num_line=20'b00011100000000000000;
                    28: num_line=20'b00011100000000000000;
                    29: num_line=20'b00011100000000000000;
                    30: num_line=20'b00011000000000000000;
                    31: num_line=20'b00011000000000000000;
                    default: num_line=20'b00000000000000000000;
                endcase
            end
            4'b1000: begin
                case (y)
                     0: num_line=20'b00000000000000000000;
                     1: num_line=20'b00000000000000000000;
                     2: num_line=20'b00000000000000000000;
                     3: num_line=20'b00000000000000000000;
                     4: num_line=20'b00000000000000000000;
                     5: num_line=20'b00000000000000000000;
                     6: num_line=20'b00000000000000000000;
                     7: num_line=20'b00000000000000000000;
                     8: num_line=20'b00000000000000000000;
                     9: num_line=20'b00011110000000000000;
                    10: num_line=20'b00011110000000000000;
                    11: num_line=20'b00111111000000000000;
                    12: num_line=20'b01111111100000000000;
                    13: num_line=20'b01111111100000000000;
                    14: num_line=20'b01110011100000000000;
                    15: num_line=20'b01110011100000000000;
                    16: num_line=20'b01110011100000000000;
                    17: num_line=20'b01111111100000000000;
                    18: num_line=20'b01111111100000000000;
                    19: num_line=20'b01111111100000000000;
                    20: num_line=20'b01111111000000000000;
                    21: num_line=20'b00111111100000000000;
                    22: num_line=20'b01111111100000000000;
                    23: num_line=20'b01111111100000000000;
                    24: num_line=20'b01111111100000000000;
                    25: num_line=20'b01110011100000000000;
                    26: num_line=20'b01100001100000000000;
                    27: num_line=20'b01110011100000000000;
                    28: num_line=20'b01111111100000000000;
                    29: num_line=20'b01111111100000000000;
                    30: num_line=20'b01111111100000000000;
                    31: num_line=20'b00111111000000000000;
                    default: num_line=20'b00000000000000000000;
                endcase
            end
            4'b1001: begin
                case (y)
                     0: num_line=20'b00000000000000000000;
                     1: num_line=20'b00000000000000000000;
                     2: num_line=20'b00000000000000000000;
                     3: num_line=20'b00000000000000000000;
                     4: num_line=20'b00000000000000000000;
                     5: num_line=20'b00000000000000000000;
                     6: num_line=20'b00000000000000000000;
                     7: num_line=20'b00000000000000000000;
                     8: num_line=20'b00000000000000000000;
                     9: num_line=20'b00011100000000000000;
                    10: num_line=20'b00011100000000000000;
                    11: num_line=20'b01111111000000000000;
                    12: num_line=20'b01111111000000000000;
                    13: num_line=20'b01111111000000000000;
                    14: num_line=20'b11110111100000000000;
                    15: num_line=20'b11100011100000000000;
                    16: num_line=20'b11100011100000000000;
                    17: num_line=20'b11100011100000000000;
                    18: num_line=20'b11100011100000000000;
                    19: num_line=20'b11110011100000000000;
                    20: num_line=20'b11111111100000000000;
                    21: num_line=20'b11111111100000000000;
                    22: num_line=20'b01111111100000000000;
                    23: num_line=20'b01111111100000000000;
                    24: num_line=20'b00111111100000000000;
                    25: num_line=20'b00000111100000000000;
                    26: num_line=20'b00000111000000000000;
                    27: num_line=20'b00001111000000000000;
                    28: num_line=20'b00111110000000000000;
                    29: num_line=20'b00111110000000000000;
                    30: num_line=20'b01111100000000000000;
                    31: num_line=20'b01111000000000000000;
                    default: num_line=20'b00000000000000000000;
                endcase
            end
            default: num_line=20'b00000000000000000000;
        endcase
    end
    always @(*) begin
        has_color = num_line[x];
    end
endmodule